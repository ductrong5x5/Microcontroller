library IEEE; 
use IEEE.STD_LOGIC_1164.ALL;


entity Project1_OR_GATE is
port --- put input and out put here
(
INPUT_A, INPUT_B : IN STD_LOGIC;
OUTPUT : OUT STD_LOGIC
);

end Project1_OR_GATE;
Architecture behavioral of Project1_OR_GATE is
begin

OUTPUT<= INPUT_A OR INPUT_B;


end behavioral;